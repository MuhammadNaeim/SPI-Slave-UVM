package shared_pkg;
    int correct, error;
endpackage
